module Xor(input A, B, output Z);
  assign Z = A ^ B;
endmodule