module Not(input A, output Z);
  assign Z = ~A;
endmodule