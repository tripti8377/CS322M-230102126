module And(input A, B, output Z);
  assign Z = A & B;
endmodule